LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom395 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom395 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom395 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"01001000",
"10101110",
"01010010",
"11100000",
"10000101",
"11100001",
"01011111",
"11100010",
"00000110",
"00000010",
"10110100",
"00111001",
"10000110",
"11011010",
"01111101",
"11001100",
"00000111",
"10111101",
"11010001",
"10100110",
"01110111",
"01010101",
"10001000",
"10110000",
"01001110",
"11100011",
"00110101",
"01111011",
"10111111",
"10111100",
"11001000",
"00010001",
"00010000",
"10001110",
"01010001",
"01001011",
"00001100",
"01101011",
"00111010",
"00011110",
"10000001",
"00010101",
"11001101",
"11011011",
"01111000",
"00000001",
"10010110",
"11110011",
"00101110",
"11111001",
"11110101",
"00101001",
"10000111",
"01101100",
"11101100",
"01110001",
"01101111",
"01110010",
"00001101",
"00110110",
"10001100",
"00100000",
"10110110",
"01100101",
"11111110",
"00100001",
"01111110",
"00100100",
"00110001",
"01010000",
"11011110",
"11010101",
"11010011",
"10010010",
"11010100",
"10010011",
"01100111",
"00100101",
"11001111",
"01101000",
"11011101",
"00010011",
"00010010",
"11101010",
"01011000",
"00100010",
"10010000",
"01100110",
"00111111",
"11001011",
"11101110",
"10111001",
"11110110",
"10011101",
"00111101",
"00010111",
"10001111",
"10110010",
"01100001",
"11000111",
"10001010",
"11110010",
"00101000",
"10100011",
"01000110",
"00001010",
"10110101",
"00100111",
"01000000",
"10000100",
"10100100",
"01111010",
"01101010",
"10101111",
"11000001",
"01000011",
"11101011",
"11110100",
"01010100",
"11111100",
"01101101",
"10110111",
"00110000",
"01110110",
"11000010",
"01110100",
"10001001",
"01101110",
"11000100",
"00000100",
"10101101",
"01111001",
"01000010",
"01010111",
"01001001",
"01000001",
"01100100",
"00010110",
"01001010",
"11010000",
"01011110",
"00010100",
"00011001",
"10111010",
"10011100",
"01010011",
"00111011",
"11011000",
"10011011",
"11111101",
"00011100",
"11010110",
"00011011",
"11010010",
"11000101",
"11011001",
"11100100",
"01000100",
"10010001",
"10111110",
"11100110",
"01001111",
"10011000",
"00101100",
"11111111",
"00011111",
"01111111",
"00101011",
"00000011",
"11111010",
"01011010",
"11011111",
"11000011",
"00111000",
"10011010",
"00111110",
"01000101",
"10010100",
"11101001",
"11110000",
"00110111",
"10100000",
"10100101",
"00011101",
"10101010",
"11011100",
"10101001",
"10111011",
"10111000",
"11111011",
"11101000",
"01100000",
"01011001",
"10011110",
"10110001",
"01011101",
"00101111",
"00101101",
"01100010",
"10001101",
"10010101",
"00011010",
"10010111",
"01110101",
"00001111",
"10100001",
"11000110",
"10011001",
"10100111",
"01011011",
"11110001",
"11001110",
"01110011",
"00110011",
"00001000",
"01000111",
"11100101",
"11001001",
"01010110",
"00001011",
"00110100",
"11110111",
"10000000",
"00001110",
"11101111",
"10000010",
"11100111",
"00100110",
"00000101",
"11101101",
"00110010",
"01101001",
"11010111",
"10011111",
"10000011",
"00111100",
"10101000",
"01110000",
"11111000",
"10101011",
"10101100",
"10100010",
"11000000",
"10001011",
"00001001",
"00101010",
"11001010",
"01011100",
"01001101",
"00000000",
"10110011",
"00011000",
"01001100",
"00100011"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;