
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY Inv_SBox369 IS
   PORT( 
      invsboxip : IN     std_logic_vector (0 TO 7);
      invsboxop : OUT    std_logic_vector (0 TO 7);
      clk       : IN     std_logic
   );


END Inv_SBox369 ;

ARCHITECTURE rtl OF Inv_SBox369 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"10011111",
"10111010",
"00100110",
"11011010",
"11000110",
"00101010",
"00000010",
"10110110",
"11000001",
"01111001",
"00010100",
"10110000",
"00100010",
"00001100",
"10111111",
"01101010",
"10101000",
"01100001",
"00110001",
"10001100",
"10100111",
"11001101",
"10011001",
"01011110",
"10010011",
"11010001",
"10111101",
"01101100",
"11011011",
"11111001",
"01111100",
"01011100",
"11110000",
"01101000",
"10101110",
"10110111",
"01111011",
"10101100",
"10010111",
"01111101",
"10000010",
"00110011",
"11110110",
"01011111",
"10010100",
"10111011",
"01011001",
"10110010",
"00100001",
"01100010",
"01001110",
"01011010",
"01010111",
"00001011",
"11100011",
"01001001",
"01001111",
"01001100",
"00001000",
"01110001",
"11110011",
"00101000",
"10000110",
"10010110",
"11110001",
"01110110",
"11010000",
"00011111",
"01100000",
"00111000",
"01100110",
"10111110",
"11010101",
"01000111",
"11000100",
"10110100",
"11010110",
"10110001",
"10011000",
"11100010",
"01010100",
"00011101",
"10001000",
"01110011",
"00011000",
"11010100",
"11111111",
"01010001",
"11101011",
"10111100",
"11011110",
"11101010",
"10000011",
"10111000",
"00100101",
"01001101",
"11110101",
"00110111",
"01101110",
"00000000",
"00001010",
"01100111",
"01011000",
"10101111",
"01111111",
"00101100",
"00011010",
"11101111",
"11100111",
"01010010",
"00110101",
"01100101",
"01110000",
"00001101",
"00010010",
"11001111",
"00010011",
"10110101",
"01101101",
"00100011",
"11011001",
"10100010",
"00101011",
"10001010",
"00000001",
"10011010",
"01011011",
"00111001",
"10110011",
"10100000",
"00011011",
"01000110",
"10101101",
"00001110",
"01000101",
"01110010",
"11010111",
"11110100",
"11001110",
"00101111",
"10010101",
"11111100",
"10100100",
"11001010",
"00111010",
"11100110",
"00010111",
"00110110",
"00001001",
"10100101",
"11011111",
"11101101",
"11101100",
"00111110",
"01110100",
"00101110",
"10001110",
"00011001",
"10101001",
"11101000",
"10000111",
"10001101",
"00010110",
"10010010",
"11100001",
"11110111",
"01010000",
"01011101",
"11001011",
"01100100",
"00101001",
"11111010",
"11101110",
"01100011",
"00000111",
"00010101",
"11000010",
"01101001",
"10100011",
"01010011",
"11010011",
"11011000",
"01111010",
"10000100",
"00000101",
"11000101",
"10001011",
"00111100",
"11110010",
"00010001",
"01111110",
"00000110",
"11101001",
"00100111",
"10010001",
"00101101",
"01101111",
"10111001",
"01110101",
"10011101",
"00111101",
"11001001",
"01000010",
"10011100",
"10101010",
"01001000",
"10011110",
"00010000",
"11111101",
"00000100",
"00011110",
"10000000",
"01000100",
"00001111",
"10000001",
"01000000",
"00111111",
"01000011",
"00000011",
"01001011",
"11000111",
"11111000",
"10010000",
"00100000",
"11010010",
"10100110",
"10011011",
"11011100",
"11111011",
"01111000",
"11111110",
"00110100",
"01101011",
"01010101",
"11100000",
"00100100",
"11001000",
"10000101",
"11000011",
"01010110",
"11000000",
"11001100",
"00111011",
"10101011",
"11011101",
"01000001",
"00110010",
"10100001",
"00110000",
"10001111",
"00011100",
"11100100",
"01110111",
"01001010",
"10001001",
"11100101"
);				  
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(invsboxip));
	invsboxop <= rom(addr_int);
  end if;
end process;
END rtl;

