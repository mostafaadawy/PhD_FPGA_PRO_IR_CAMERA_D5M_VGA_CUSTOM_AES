LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom357 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom357 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom357 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"11000000",
"01011110",
"10110010",
"01000000",
"11111101",
"01011010",
"10100111",
"01110100",
"11011110",
"10111011",
"00101100",
"11010110",
"11010011",
"10110101",
"00000001",
"00011001",
"11000100",
"11100000",
"10010001",
"11011101",
"00100011",
"00111000",
"11101000",
"10110110",
"10010101",
"01101110",
"00111011",
"11010100",
"00001000",
"11101101",
"01111110",
"11100110",
"01110010",
"10011010",
"10011100",
"01010001",
"10001110",
"11110001",
"00011010",
"10001100",
"00010000",
"00011000",
"01000011",
"10101111",
"11001110",
"10000110",
"10001010",
"01001011",
"10001001",
"10000010",
"00110100",
"00101010",
"11001001",
"11100111",
"01001111",
"10011101",
"10010100",
"10011000",
"11111010",
"00111101",
"00100100",
"00001001",
"11000001",
"10111010",
"10100001",
"01101101",
"11101011",
"10000001",
"10011111",
"01100001",
"10110000",
"00000100",
"01010110",
"11111110",
"10111001",
"00000010",
"00000110",
"10010010",
"11110011",
"00101101",
"10111000",
"10000100",
"11110110",
"11000011",
"11110010",
"00101000",
"01011111",
"00011111",
"00000101",
"01100111",
"10011001",
"00111010",
"10111101",
"01101100",
"10010111",
"00101111",
"01011011",
"11010111",
"00010110",
"11001011",
"10010011",
"01111000",
"11100100",
"11011010",
"11000111",
"11110100",
"00110110",
"11101001",
"00100001",
"01000101",
"01110101",
"11110111",
"00110000",
"01000111",
"10110100",
"01111011",
"10011110",
"11011000",
"10000011",
"11100011",
"01100000",
"00001110",
"11101100",
"01001010",
"01111010",
"00111001",
"00110010",
"01010101",
"10100011",
"01010010",
"00101110",
"01110111",
"01001000",
"01001100",
"00001011",
"00010100",
"00010010",
"00101011",
"00110001",
"10001111",
"01100010",
"11100001",
"10100110",
"00111111",
"11010000",
"00100111",
"11111001",
"10000000",
"10101101",
"00000000",
"00100010",
"11110101",
"11111111",
"10101100",
"11010001",
"00100101",
"10011011",
"01101011",
"00000111",
"01000110",
"01101000",
"10010000",
"10100010",
"11110000",
"10111100",
"11001101",
"10101001",
"01101010",
"00110011",
"11111000",
"10000111",
"10110111",
"11000110",
"11001100",
"01111101",
"01001001",
"01011101",
"01000001",
"01010000",
"10010110",
"01001101",
"11010010",
"00011110",
"10001101",
"11001111",
"00111100",
"00001100",
"00100110",
"11001000",
"01111001",
"00110101",
"00001101",
"01101001",
"00011100",
"01010011",
"10101110",
"00010101",
"00000011",
"11011001",
"10101010",
"00110111",
"00010111",
"00011011",
"01011100",
"11101110",
"11000010",
"10100000",
"11111011",
"10111111",
"11000101",
"00011101",
"00100000",
"10101000",
"10001011",
"11100101",
"11101010",
"00001010",
"01110110",
"01000010",
"11011111",
"01110000",
"00010001",
"01000100",
"01100110",
"00101001",
"11011100",
"11001010",
"01100100",
"01110001",
"01010100",
"10001000",
"01011000",
"01101111",
"01111111",
"10110001",
"01010111",
"10111110",
"10000101",
"00010011",
"01100101",
"00001111",
"01011001",
"11100010",
"00111110",
"11010101",
"10101011",
"10100100",
"10100101",
"11011011",
"10110011",
"11101111",
"01110011",
"01001110",
"11111100"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
