LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom375 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom375 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom375 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"00100111",
"11100100",
"10001010",
"00011110",
"10100000",
"11011110",
"10010111",
"00001000",
"11011101",
"10111110",
"01001001",
"00000111",
"01110110",
"10110111",
"11010010",
"11010000",
"00011101",
"11100110",
"11110111",
"00001111",
"10001101",
"11001101",
"10111101",
"10001100",
"01010001",
"11001000",
"00100010",
"00101000",
"00001001",
"00111101",
"10111011",
"11011011",
"10111010",
"11000010",
"01011100",
"00010001",
"10100001",
"10100101",
"00101001",
"11111010",
"01010101",
"10110100",
"11011111",
"01110111",
"11111111",
"01010010",
"00001100",
"01000101",
"01011111",
"01111111",
"10110001",
"01101101",
"10110110",
"11100001",
"11000011",
"10001011",
"11000110",
"01101001",
"10011101",
"01010111",
"10000111",
"01000111",
"11000100",
"10000000",
"00111111",
"11010110",
"01000100",
"10101010",
"10110011",
"00000010",
"11111100",
"00001110",
"10010001",
"00111011",
"11001001",
"10011010",
"00000000",
"10010101",
"01000110",
"10101011",
"01100100",
"11110011",
"01111000",
"11100101",
"10001000",
"10000100",
"11110110",
"11100010",
"10100010",
"01110101",
"00101101",
"11000101",
"00110000",
"00010100",
"11010100",
"10011000",
"01110000",
"11110100",
"01111101",
"10001110",
"10100110",
"01100001",
"11000001",
"00100001",
"10101111",
"00010101",
"10001001",
"10010100",
"11101001",
"10110010",
"00110011",
"11111110",
"00010111",
"10011011",
"01111010",
"00100011",
"01100110",
"01101111",
"11010111",
"01010100",
"01111001",
"11101011",
"11011010",
"11010001",
"01110001",
"01011010",
"01111011",
"01110100",
"10010010",
"11001111",
"10000110",
"00000110",
"01110010",
"00001101",
"11110000",
"00101111",
"01001100",
"00000011",
"11000000",
"00011011",
"00011000",
"11100111",
"10101100",
"11111001",
"11010101",
"01100101",
"00011010",
"10111001",
"01001111",
"01100000",
"00110110",
"01100111",
"10011111",
"10100100",
"00011001",
"10010000",
"11010011",
"00101110",
"11110001",
"11101000",
"11001100",
"10111000",
"00101011",
"10011100",
"11100000",
"00100101",
"11101110",
"00010000",
"00100000",
"10000101",
"10010110",
"11011100",
"01011011",
"11000111",
"10101001",
"00101100",
"01101000",
"00000100",
"01001000",
"11110101",
"10100011",
"10111100",
"10001111",
"10011001",
"11111011",
"01011101",
"11001010",
"00111100",
"11011000",
"10110101",
"01110011",
"10000011",
"10011110",
"10110000",
"11101010",
"10000010",
"10101000",
"11011001",
"10100111",
"00110001",
"01011110",
"00111001",
"10000001",
"00001010",
"01100010",
"00100100",
"00110010",
"11001110",
"01000010",
"00111000",
"00000101",
"01111110",
"01011000",
"11001011",
"00010110",
"00110111",
"01010011",
"00110101",
"11101101",
"00100110",
"01000000",
"01010000",
"01001011",
"01001110",
"10101101",
"11111101",
"01011001",
"01001010",
"00011111",
"00000001",
"11101111",
"00001011",
"01000011",
"11100011",
"00101010",
"00011100",
"10101110",
"00010010",
"11110010",
"01000001",
"11111000",
"01010110",
"01101110",
"00010011",
"11101100",
"01101011",
"10111111",
"00111110",
"00111010",
"01001101",
"01101010",
"10010011",
"00110100",
"01101100"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
