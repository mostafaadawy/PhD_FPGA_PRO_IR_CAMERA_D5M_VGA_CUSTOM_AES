LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom397 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom397 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom397 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"01101001",
"10010000",
"01100110",
"00110010",
"10011010",
"00001110",
"01100100",
"01000001",
"11001011",
"10101001",
"10011111",
"11111010",
"11010101",
"10101010",
"01100101",
"00100100",
"11110111",
"01110111",
"00110111",
"00011101",
"10000011",
"11101011",
"10011000",
"00011010",
"00101010",
"01111101",
"10111101",
"00100101",
"00000010",
"11101110",
"11100101",
"11100111",
"01000101",
"01010000",
"00101001",
"11000100",
"11101100",
"10100111",
"11001100",
"11110000",
"01011100",
"01001101",
"00010011",
"10010110",
"10100010",
"00001001",
"10011110",
"11111111",
"01011010",
"10100001",
"11000111",
"01101111",
"11101001",
"00010101",
"00001100",
"00011011",
"11000101",
"10010111",
"01010110",
"00010100",
"10100101",
"10110110",
"00100000",
"11010110",
"00100001",
"00010001",
"01110000",
"00001101",
"01111111",
"01001110",
"01000110",
"01010010",
"00110101",
"01001011",
"10100100",
"11001001",
"00000001",
"00011110",
"00110001",
"00001111",
"00101111",
"00010111",
"11111100",
"11011011",
"01110100",
"00110000",
"11011110",
"01001000",
"00011100",
"10010101",
"00000110",
"01010011",
"11010011",
"01100111",
"00011000",
"11111101",
"00101101",
"00011111",
"01111010",
"10001101",
"10000111",
"01110101",
"10110100",
"00100110",
"11100000",
"01110001",
"10100011",
"10000010",
"01011000",
"00000111",
"11010100",
"10111010",
"11011010",
"10101000",
"10110101",
"11011001",
"10011100",
"11001111",
"11111001",
"01100000",
"11011000",
"00010010",
"00000000",
"01111001",
"10001001",
"00000100",
"11000010",
"10111000",
"00111100",
"01100001",
"01000010",
"01110110",
"11011111",
"01101100",
"11101010",
"01001001",
"01010100",
"01100010",
"11101000",
"10110011",
"11110101",
"00001011",
"11110001",
"00101000",
"01111110",
"11010010",
"11001101",
"00100011",
"11110010",
"10001110",
"10000000",
"11111000",
"00110110",
"11100011",
"11010111",
"00100010",
"11011101",
"11110011",
"01001010",
"00101110",
"01010101",
"00010000",
"11000000",
"10110001",
"01011001",
"01000011",
"10101100",
"01101000",
"00111111",
"10111011",
"01101101",
"10101111",
"11001010",
"11000110",
"00111000",
"10111001",
"01110011",
"10101110",
"11011100",
"10111100",
"10011101",
"11000011",
"11010001",
"01001100",
"11111110",
"10100110",
"00111011",
"10010010",
"11100100",
"00101011",
"01011011",
"11111011",
"00101100",
"11110110",
"11000001",
"10110010",
"01011101",
"10001111",
"11101111",
"01111000",
"10010001",
"01011111",
"10010100",
"01110010",
"11101101",
"01000000",
"10001000",
"10110111",
"01000100",
"00110100",
"00100111",
"11100001",
"01101010",
"00000101",
"10000110",
"11001000",
"10010011",
"10001010",
"01111011",
"10000100",
"01010001",
"11100110",
"00111101",
"10011001",
"00001010",
"00110011",
"10111111",
"00111001",
"00000011",
"10001100",
"00001000",
"01101011",
"00111110",
"10000101",
"00011001",
"11001110",
"10110000",
"10001011",
"10101011",
"10100000",
"11100010",
"01000111",
"10111110",
"01001111",
"01011110",
"10011011",
"01010111",
"10101101",
"01101110",
"10000001",
"00010110",
"00111010",
"11010000",
"11110100"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;