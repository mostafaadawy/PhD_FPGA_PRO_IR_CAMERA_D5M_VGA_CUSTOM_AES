LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom355 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom355 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom355 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"11100001",
"01100000",
"00101111",
"01100010",
"11100010",
"01101000",
"01001000",
"01101100",
"11100011",
"00110100",
"10101110",
"00101001",
"11100110",
"10010101",
"11111011",
"11001110",
"11101001",
"10001111",
"00101110",
"00001101",
"11000101",
"01010011",
"10000101",
"01001101",
"01000110",
"01100110",
"10100001",
"10100111",
"00010101",
"11101011",
"00100010",
"00011011",
"10111000",
"00010110",
"00101011",
"10100101",
"00011000",
"11010110",
"11001000",
"10011101",
"01010100",
"01111001",
"00111101",
"10011111",
"01110110",
"01100101",
"00011101",
"00010111",
"01110100",
"00001110",
"11110001",
"00110001",
"11101100",
"01010001",
"00001111",
"10001100",
"00000001",
"10101011",
"01011000",
"01000011",
"00101010",
"10110000",
"11000011",
"11011011",
"01010010",
"01101010",
"10000011",
"00110010",
"11011001",
"10001010",
"01000111",
"11101010",
"00000000",
"00110000",
"11010011",
"11010010",
"10110100",
"10110111",
"10110110",
"10000001",
"00010001",
"01001111",
"11111000",
"10110001",
"01101110",
"00000010",
"01000001",
"01111011",
"00010000",
"10010110",
"11100100",
"10001101",
"01101101",
"01011011",
"01011100",
"11110101",
"01011001",
"01001011",
"11100101",
"10111001",
"11010101",
"01000000",
"00100111",
"00000110",
"01001010",
"10101001",
"10100100",
"11000100",
"01110111",
"00100001",
"01010101",
"10011110",
"10011001",
"01010110",
"01011111",
"00000101",
"00001010",
"00110111",
"11110011",
"00101100",
"01111110",
"11000000",
"11000111",
"10011100",
"10000111",
"00010100",
"00110011",
"01001110",
"00111111",
"11001100",
"11110110",
"10110011",
"11100111",
"00110110",
"00010011",
"10011000",
"11001011",
"10101111",
"00111110",
"11111101",
"10010111",
"10000110",
"01110001",
"00001000",
"10101010",
"11000001",
"11011111",
"01110000",
"11001010",
"00011010",
"00111011",
"10100110",
"10111011",
"11011100",
"10001000",
"01001001",
"00001001",
"10111110",
"10001001",
"10010011",
"00010010",
"11101110",
"01010111",
"10000100",
"01110101",
"10011010",
"10100011",
"10001011",
"00000111",
"11011101",
"11101000",
"10111100",
"11011110",
"00100011",
"01111111",
"01011101",
"01101111",
"01100001",
"11010111",
"01100111",
"10010100",
"11110111",
"10100000",
"00111000",
"00011001",
"10111111",
"01101001",
"00100101",
"01110010",
"11110000",
"11111100",
"10111010",
"00101000",
"11110100",
"01110011",
"10011011",
"01111010",
"00111010",
"00100000",
"11001101",
"00000011",
"10100010",
"00110101",
"11010100",
"11111111",
"01011010",
"01001100",
"11010000",
"11010001",
"10010010",
"11111010",
"00100100",
"00001011",
"00001100",
"10000000",
"00000100",
"10111101",
"11101101",
"01100100",
"10101101",
"01000010",
"11111110",
"01111000",
"10000010",
"10010000",
"10101100",
"00011110",
"10101000",
"11111001",
"11000110",
"01111101",
"00011111",
"01010000",
"01101011",
"11011010",
"11001111",
"01000100",
"11101111",
"00100110",
"00111001",
"11001001",
"11000010",
"11100000",
"10001110",
"10110010",
"01011110",
"00111100",
"10110101",
"10010001",
"01000101",
"00011100",
"11110010",
"11011000",
"00101101"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
