
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY gen_rom IS
port(
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 63)
	 );
END gen_rom ;

-- hds interface_end
ARCHITECTURE rtl OF gen_rom IS
 Type rom_type is array (0 to 255) of std_logic_vector(0 to 63);
constant rom : rom_type :=(
"1011110110100111001010001111010011100001001101101001010111000000",
"0011000110001101101001100101111100001011001001111001111011000100",
"1100011000101111000101011101100000110000101101000111101010011110",
"0100101111100010100000010101111101100111101011011001000000111100",
"1101111101110101000000011010100001101100001110010100101111100010",
"0101010000111011100011110001111010010000110101100010011110101100",
"1101100011111011110010010101010001110011101000001110001000010110",
"0110111010100000010110110001111111001001010011010011001010000111",
"1110001001100100110010010111100011110001001110110000101011010101",
"0110011100001001010010001111111000011011110101011100001000111010",
"1111101110101001100000110100011000011110011100101100110101010000",
"0111000010001110001100101101111101010110100100010100101011001011",
"1111010100100001101000000110100110001100001111101101101101000111",
"1000101011010100000011111011111001100001110001110101001000111001",
"0000111010001001011111000010011010110101101000110100111111010001",
"1001001101001100111110101000111010110111001000001101000101010110",
"0001100011111110011001110000100111010011001011001010101101000101",
"1001110110100010111001010111111100000110101110000011000111000100",
"0010000101101000010101111111101000111110101110010000110111000100",
"1010010100001001110100100111111101000011011010001100101100011110",
"0010101111001101001100001110011101101001000101001000111110100101",
"1011111101100000101011100100110101110001100111000010010110000011",
"0011010100100110000111011100100110110111100011101111101000000100",
"1011100011010110100110100010111111000111000101000011010100001110",
"0100110110001010000001111011011011110001111000110010110010010101",
"1100001001001110011101100001111100001001101111011010010100111000",
"0100011111110001111001011001100000101101011010111010110000000011",
"1101101110000100010100010000111101100011011110100010110011101001",
"0101000001101001111000011000101001111100111100111101001010110100",
"1110010000001011010111011100111101111010011000011000001100101001",
"0110101011001111101110010011010110000010010011100001000011010111",
"1110110101100010001110101011111110010111000010001100010001010001",
"0111001100011000101110010100101011110000111001101100001001011101",
"1111011111001000000101011010111000000110100100110100101100101101",
"0111110010001101011000100001100100111110010100000100101011111011",
"0000001001010001001101101011010010011000011111101101111110101100",
"1000010111110011011100000001101010011011110101100100001011001110",
"0000101110010110111011010101000110001111011100110010110010100100",
"1001111101001010010111001110011010000010000100001101001110110111",
"0001010000001110110010100110001011011001001111110111101101011000",
"1001100011000001010001111110011011110000101110100010001111010101",
"0010110101100101101101110011000000011001101011001111111010000100",
"1010001000011000010001011101100100111110011001111100000010111111",
"0011011111011011100100010010000001100100111101011000111010101100",
"1011101001111111000000011001011001011000110111101100001101000010",
"0011000001010100101011100001001010111111100010011100110101100111",
"1100010011100101111110100111011010010001001000111000101100001101",
"0100101010011000011010111111000011010111111000011100010100110010",
"1100111001001011110101100101011111111010001110010010000110000000",
"0101001000000001011110011110001101001010101111011000111101101100",
"1101011110110010110000110101100000011010000010010100111011110110",
"0101110001100111001000011101000010000011111110011011010011101010",
"1110000100101010101100000101100001111001110000110110110101001111",
"0110010111011110000111001001000010001011010011110010001101111010",
"1110100101110001101011000010011010110011000011011111010110000100",
"0111111100100100000010101001000111011000110001100101001110111110",
"1111001111010111011010001110010111001011010000000001100100101010",
"1000100110101100111101000101000000010110001111101101001010110111",
"0000110101011111011000111100100000101010000110111001011111100100",
"1000000100000011111001000111001010010101110110110110101011001111",
"0001011110110101010011111100100001100011100100101110110110100000",
"1001101101011000110011100010000001111101001100011010010011110110",
"0001000000111101010111001010100010110010111111100110100101000111",
"1010010011010000100110000010000111100111110010111111001101010110",
"0010100110000011000110101011011111111110010101101100110101000000",
"1010111000100110100001000000000100110111100110111100010111011111",
"0011001011101010000001011000100101001100111111010001101101100111",
"1011011110011110010100011111000001001101100010100110001011000011",
"0100110001010000111011110110100101110011100010100010110110110001",
"1100000011110100011011011011000110001010001001010011100101111110",
"0100011010111000110111000010100110100000111100011110011101010011",
"1101100101011011001110001100000011100110011111110010010010100001",
"0101111100011110101001110010100111011011010010000000110000110110",
"1101001111000001001001101010000001000111010110111111100110001110",
"0110100001110100101100100000110000111010111001011101111110010001",
"1110110000101000000000111001000101101111101001000101101101111101",
"0110000111101100100011111101011101000011001010111010000001011001",
"1111011010011110110110110100000001111000000101011010001111000010",
"0111101101000010100011001110100110100000110100110101000111110110",
"1111111011010101101101110011000010100100011000011100100000101001",
"1000010010111010001101111101100111101100000111110101000001100010",
"0000100101101110110001000010000111110011110110100111100010110101",
"1001111000010000010001011011101000101000110101110011011011001111",
"0001001111000101101100100000010001111111100110001101101001101110",
"1001011001111000000111111010101100110010010000001100010111101101",
"0010110000111011100011101111000001101001110110100001011101000101",
"1010000011101101000110010110100001111111010110111100001000110100",
"0010011010100001100010111110000011000101011101001001111111010011",
"1011100100110101111101110100101011011100000000010010011011101000",
"0011111011111000010101001011000011010001110010101001011100100110",
"1011001110101100111000100100100000000111100111010110000111110101",
"0100100001101111001100001011000101011101100110100010111011000111",
"1100110100010011101011110010100001010100000001111110011010011011",
"0100000111000111001111101001000010001010110100101011111101010110",
"1101010101111010100110110000100001101111010011100010001111000001",
"0101101100101101000110010111000011000110010011101111101000111000",
"1110111111000000011101011101100010100110000101001001001100101011",
"0110010010010011000001111000000111110010110101011011111011001010",
"1110100000110111011000101101101000000101100111110001101111000100",
"0111110111111001110000000011000101001011010110101000111000100110",
"1111001010101101010111101001011100110001110001100100100010110000",
"0111011001010001110111100010001110011010110001000000100011111011",
"0000110000010110010110111010100110001111010000101110011100111101",
"1000000011001001101101110001001111010100010111110110001010101110",
"0000010110001100001001111010101111101001111101100001010011010011",
"1001101000101111100001001110000111011100011001011011000000110111",
"0001111011010011000001011000101000100111100101101100101101001111",
"1010001110000110100100001110001001001101000101010111101111111100",
"0010100001001010111111100011100101010000110110111100011001110001",
"1010110011111011010110011000000101000110011100111101000000101110",
"0011000110110000111010100100100110001101010101100111111111000010",
"1011010101000011011010101100000111010010000001111111100011101001",
"0011101100001000110101100001101011101001110011110101011100100100",
"1100111110101000001001000111000111101101011010010011000001011011",
"0100010110001110101100101111100100000110001110100001110111000111",
"1100100000100001001100001001010101101101010010101110011110111111",
"0101110111000100100011111011011100100000101000010110111000111001",
"1101001010000111000011000101001110010110101011110001101111100100",
"0101011100111100100010111101100101101110000101001111101000100000",
"1110101111111101110001100010000110000011101001000101011100001001",
"0110000010110011011110001100101011100101110100010010111110010100",
"1111010001010111110100110001001011101100100010111010011010010000",
"0111101000001001010000101011110000010101011011101101111100111000",
"1111110110101011100000000001001101001001111001100010011101011100",
"1000001101110000010011111001101101011110101000101101110001100001",
"0000100000100101101111011111001101110110100100011100101001001110",
"1000110011010101000110100100100101111110000011110011001001101011",
"0001001010011011100001111110001111000000111110101101010101100100",
"1001010100111110111101100010101011000111100000011011000011010100",
"0001101111110010011101011100001111101010010000001000100101101101",
"1010111110000011110100010010100100000101010011100110011111001011",
"0010010001101001011100001100001101011101111010111010100011110001",
"1010100000001100110111110001011101001110011001010011001010011011",
"0011110110111111010010100110000101110101001010000000110010011110",
"1011001001110011110010101111100101101000000000011110010011010101",
"0100011100010110001010101000001111010000111011111001110001011011",
"1100101011010111100001001110100110110010001101100000000101011111",
"0100000010011101000101100101001111111100011110101110101110000010",
"1101010000110000100100101100101100010110111101111010010111101000",
"0101101011100010111100000011010001101001110011010001101101111000",
"1101111010000101010011001001101000101111001101111011000001100001",
"0110001001011011111011000000001110000100011110101101111110010001",
"1110011100001101010010101000101101101001111100100011010100011100",
"0110110010110001110101111111001010010000100000111110101001000101",
"1111000101100100001110001001110011010101011111101010001010110000",
"0111010100011001110001001110001011111011000010100110110100111000",
"0000101011011011001000110110110000010100111110000101100101111110",
"1000111101111110011000001011001000111001101001001100110101010001",
"0000010001010010000111100111110010001101011000111010101111111001",
"1001100011100100011011001010000101010010000011010011111101111011",
"0001110110011000111110100010101101100111110001001110001101010000",
"1001000101011101011010001010001011001111011100110100000011101011",
"0010011100000001110110000011110011100110010101001001101110101111",
"1010101110010010010000110111000111111100000011101101010101101000",
"0010000001111000110000111111101100010100110110101001011011100101",
"1011010000011010001100000111010101101100100111010010100011101111",
"0011100111011110100011001011011100101010000101001111010100000110",
"1011111001110000001011000100001110000101111100011010011011011001",
"0100001000110110101010111100110110000111111011110000100101010001",
"1100011111100110111101010001001010101101010010011011000000111000",
"0101110010011011011001001000110111100001001000111010111101110000",
"1101000001011110110000110001010011111001101100100111011010101000",
"0101011000000010100000111010110100010100110011111110101101111001",
"1110100110100100110000001111001000110110011110111000000101011101",
"0110111101011001001011010100101100111100000010000111111010100001",
"1110001100011100101010111101001001100000111101010100011110001001",
"0111100011011111000110010011101101100101101000001100111000100100",
"1111110001100010100101111011001110101101000111100100010110000000",
"0111000100111000000010010100110111100101001011000110111110111010",
"0000011111101010100000111011010011111001110001011101001000010110",
"1000101110011101111100010000101000101110011000110101110001110100",
"0000111101010001011111101001010000111000011011010010101111001010",
"1001010011110011110111001110100000100111000010101011011000010101",
"0001100110110111010011010110001110000000111010101100010100101111",
"1010111001011011110001111101100001000011001000010000111110010110",
"0010001100011110010110010111011011001101010000001111101010001011",
"1010011011010001101101011100100111100010111110000100000000110111",
"0011110001110101000101000110100011111010110110110010100111100000",
"1011000000111001100000101100110111111110010101101010000101110100",
"0011011011101011000011110010010100010111100010011100101001001101",
"1100100110001111010111010110101000010111111010110010000001000011",
"0100111000110010111110110000011001110001101011000101100111011000",
"1100001111110110010110010111101101000010100010101101000000011110",
"0101100010111010110101101111001001111100000000110100111000011001",
"1101110001011011001101000110101010010000111100010010011111101000",
"0101000100100000110001101101011111101001101011111011100000110100",
"1110010110110011001000010110110011111101010010010111000010001010",
"0110101101111000101011111001001000000011000111000100111011010101",
"1111111000101001000111000011101001001000101101011101000001110110",
"0111010011101101100010100110001000111111100100001011110000010101",
"1111100010010001111001110000101101010100001111010010011011001010",
"1000110100110101011110010110001010111100000010101111111001000001",
"0000001111111001110101011110101010000001101101000111011000101100",
"1000011010111100010000100101001111101001011100001010111100011101",
"0001110001101111101100101101100111101000001110100111010001010000",
"1001000000010100010111110110011100101000111011001011110100111010",
"0001010111000111101111101010100100100110110101000011100000001111",
"1010100101101000000111000010010001011111011100110000111011011011",
"0010111000111100100110001010101101010100000000011101011111110110",
"1011001111100000000110000010011010101100111111010101010001111001",
"0011100010010100101001011011111011000000011111010001011011110010",
"1011110000110110111100101110010010100101011100011101000010011000",
"0100000111111010011000001000110111101011001000110111100101011100",
"1100010110101110110111111001001000000001101110000011010001100111",
"0100101101100001010111100111110100101001101011001111001110000000",
"1101111100000101101110011010001101001110001001111000000101101100",
"0101001111001000001010100100111001110001000010010110110110111111",
"1101100001101011100101011010001001111100111000001111000101000011",
"0110110100101111000101010011110010101110100010110111100101000000",
"1110001011000011100001001001010111010110000110110111000010101111",
"0110011110010100000000011111110111101010001010001100101101010011",
"1111101000111000011011100101001000000001110001001011011111011001",
"0111000011111100111010111010100100100101010011010011100000010110",
"0000010110110001011111000110010010001110001111010010100110101111",
"1000101001000011110110011100111001010001111101100111101100100000",
"0000111000010111010110000100011010111010110100111001001011001111",
"1001001011001010101101001000111001111111001100000001110101010110",
"0001100001111110001101000010011011011001000011111100101010110101",
"1001110000100001101000001000111011110111110101100100101101010011",
"0010000111010101000011110011011101000110101110101000110010011110",
"1010010110000111100111010100111000010011011000101111110010110000",
"0010101001001100111110011110001101011011000000011000011111010110",
"1011111111101101010101110011101001000000110010000001100100100110",
"0011010010100010111001111101010110011000101101101111000100001100",
"1011100001000101011000110010111011001111000101111010000011011001",
"0100110100001001110000111011010111100010000101101000101001111111",
"1100000110111101001100000100111011111000100110100111001001010110",
"0101011110000000110011111010001100011110100110110110010011010010",
"1101101000010011001011000000111001010111011010011000010011111011",
"0101000011010111101010111000001101001110000101100010110010011111",
"1110010010001010000010011111110001010001101100100111001111010110",
"0110100100111110011101011000001010111010010011110001110011010000",
"1110110111110000110001001010100101111000001001010001001101101011",
"0111001010100100011000011000100111100011111101011101110000001011",
"1111011101001000110100001011110011100101100100010011001010100110",
"0111110000001011010011110010011000011110100011010011101001011001",
"0000000111001111101110101000110100110101001010011110010001100111",
"1000010101100001001111000000100101111101111110101011111001000010",
"0001101000100110101110011000111001010000110001000011011111111101",
"1001111111000111000101011110010010000011011000001101101100101010",
"0001010010011101100001010111111010111100000011110110001010100011",
"1010011100111111000000101101011011000001111010010101101110000100",
"0010110111100011011100000110110011111000100101011011010000011010",
"1010000110010110111111101011010000001101001100101000110001010111",
"0011011101011011011011010010111000010100000011111001101011001000",
"1011101000001110110010000111010000111001110101100001111100100101",
"0011111110110000010110000010110101111110100101101010010000011100",
"1100010001100011101101111001010110100010000110001101111111100000",
"0100100100011000001101100000111011001101001001010111101111111010",
"1100111010111001011100010101010011010000101011111000001000110110",
"0101001010011110000000011111110011010111011010100100100010110011",
"1101011000100001100111100101011100001100010010100011100011111011",
"0110110011100100111110101011100100010010110100111000010100000111",
"1110000010011000011010110011010101001010110111110111000100101100",
"0110010101001101111010001011110000111111001010010000011110100001",
"1111100100001110010101100010011110100100000110111101001110001100"

);

BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl; 
