LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom361 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom361 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom361 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"10000010",
"00100010",
"10010011",
"01011100",
"11000011",
"01001110",
"00011011",
"01111000",
"11111100",
"01110011",
"00110011",
"11001100",
"11110101",
"10001001",
"00110001",
"10001110",
"11101110",
"10000001",
"10101100",
"10011110",
"01101011",
"11111001",
"01001011",
"11000101",
"11011010",
"01101010",
"00101000",
"00100111",
"00010110",
"00111000",
"01001010",
"11100001",
"11111011",
"01001101",
"10100101",
"01101100",
"00010010",
"10100000",
"10000100",
"00000100",
"11110011",
"00000001",
"01100111",
"10011011",
"01000000",
"00011010",
"00011001",
"11101101",
"01011110",
"11000111",
"10111111",
"11000010",
"11100111",
"11010011",
"11000110",
"11101010",
"00101111",
"01011000",
"11011001",
"10010110",
"11001110",
"10000011",
"10011001",
"01110111",
"01001100",
"11010111",
"01000001",
"01010000",
"01110100",
"11001111",
"00000000",
"10001100",
"10001010",
"10101111",
"10110101",
"11000001",
"11101100",
"01011001",
"11111110",
"10000000",
"11010000",
"11100110",
"01000101",
"10110100",
"00111100",
"11100101",
"00001111",
"10111000",
"00011111",
"01000011",
"10011100",
"11001011",
"10110001",
"01001000",
"00110000",
"10101000",
"00100100",
"11100010",
"11111101",
"01111001",
"01011111",
"00100101",
"00001101",
"11011101",
"10110011",
"11110001",
"00100001",
"01010001",
"00111011",
"01100110",
"11011111",
"11111111",
"11001001",
"01100001",
"00101011",
"00010001",
"10010000",
"01111111",
"00111110",
"11011100",
"11110111",
"00001010",
"11011011",
"11110110",
"00010011",
"00001100",
"00011110",
"01000110",
"00000111",
"01101001",
"11110100",
"01100000",
"01010111",
"11101111",
"00011100",
"01101101",
"10010100",
"10111101",
"10000110",
"10111011",
"01011011",
"10000111",
"10111100",
"00100110",
"11111010",
"00010111",
"10010111",
"11010110",
"00000101",
"00111010",
"00001000",
"00100011",
"00110010",
"11101001",
"10100100",
"01101000",
"00010000",
"10110010",
"10101101",
"10100111",
"10010010",
"10010001",
"10111010",
"11100011",
"10100001",
"11100100",
"01110000",
"00010101",
"10001000",
"01111110",
"10100010",
"00101010",
"00100000",
"11011110",
"01010101",
"10011111",
"11100000",
"10110110",
"01011101",
"00111101",
"00011101",
"00111001",
"11110010",
"01110001",
"00110111",
"00001001",
"01100100",
"10100110",
"10011000",
"01010110",
"11001010",
"00001110",
"11101000",
"01101111",
"10101110",
"11110000",
"11001101",
"00011000",
"00101100",
"11111000",
"01101110",
"00000110",
"01111101",
"10010101",
"00101110",
"10001101",
"01010100",
"01110101",
"01010010",
"10111110",
"01100101",
"01111011",
"01000100",
"01001001",
"01000010",
"10011101",
"00010100",
"01110010",
"01001111",
"11011000",
"10001111",
"11101011",
"01010011",
"10000101",
"00101101",
"11000100",
"00110110",
"01011010",
"01100010",
"10110000",
"01000111",
"10110111",
"00110100",
"11010101",
"10011010",
"11001000",
"00000011",
"00001011",
"10100011",
"00000010",
"11010010",
"01110110",
"00101001",
"10101011",
"10111001",
"01111010",
"00111111",
"10101010",
"10101001",
"11000000",
"00110101",
"10001011",
"11010100",
"11010001"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
