LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom419 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom419 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom419 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"11000101",
"10100111",
"00011001",
"00010001",
"00000001",
"00010111",
"01110111",
"01001111",
"01110011",
"00011000",
"01111011",
"11110011",
"01011001",
"10110010",
"01000000",
"00101100",
"01110101",
"01110000",
"01101011",
"11111110",
"11110111",
"00010011",
"01101111",
"10101100",
"00000010",
"01001001",
"01010111",
"01001010",
"10100010",
"10010000",
"11011011",
"00110010",
"11101101",
"10101111",
"01000001",
"01111010",
"11101010",
"10110101",
"01100111",
"01111000",
"10101101",
"11011001",
"00101001",
"10110100",
"01110010",
"01100001",
"01001100",
"10110110",
"10000100",
"01101000",
"11111010",
"10100011",
"01011111",
"10001101",
"01111001",
"10000010",
"11011110",
"00101011",
"10101010",
"11000010",
"10011010",
"00100110",
"00111111",
"10010001",
"11001011",
"00111001",
"00100100",
"10100110",
"00000101",
"11001101",
"01011011",
"10001010",
"11101111",
"11000011",
"10001110",
"10100100",
"00001000",
"00100001",
"01001000",
"00001001",
"11101110",
"11100001",
"00000100",
"10101011",
"00111110",
"00011110",
"01000110",
"11000110",
"10001000",
"00111100",
"11101011",
"01011000",
"01100010",
"11011100",
"11110100",
"11001110",
"10001001",
"10011101",
"10111001",
"11011000",
"11100110",
"11010010",
"10000110",
"11100000",
"00101010",
"01110110",
"01111101",
"11110000",
"00111101",
"01011010",
"01101110",
"01010011",
"10010011",
"00100011",
"10010100",
"11111011",
"01000111",
"11010001",
"10101110",
"00101111",
"10110011",
"01101010",
"10011111",
"11000100",
"11101000",
"11001111",
"01100100",
"11111000",
"00011010",
"11111001",
"00110111",
"10111101",
"01001110",
"00110000",
"11101001",
"01001101",
"10000001",
"01101001",
"01010000",
"10011011",
"00011101",
"01001011",
"01010110",
"01010100",
"10010111",
"10001100",
"00100101",
"01101101",
"00110011",
"10010010",
"10111100",
"00001101",
"10000000",
"00101101",
"11111111",
"10111111",
"01000010",
"11011010",
"11011111",
"10000111",
"01111111",
"11001001",
"10100101",
"00000111",
"00001011",
"11110110",
"11010000",
"00001100",
"00101110",
"01100000",
"11100100",
"11001010",
"11011101",
"11110101",
"11110001",
"01110100",
"10011000",
"00001111",
"10010110",
"01100110",
"11100101",
"00010010",
"00001110",
"00011111",
"11010111",
"11010011",
"11100011",
"01011110",
"10010101",
"01011100",
"10101000",
"11000001",
"10011100",
"00000011",
"00010110",
"01010101",
"00110101",
"10011110",
"00100111",
"11001000",
"10111110",
"10110000",
"10100001",
"11110010",
"10111011",
"00100000",
"10111000",
"01011101",
"10001011",
"11010101",
"11000111",
"00111011",
"11000000",
"00010000",
"01000101",
"11111101",
"10000011",
"00001010",
"01100101",
"11111100",
"11010110",
"00110001",
"11001100",
"00111000",
"01010010",
"00010100",
"00011011",
"00110110",
"01000011",
"01000100",
"10110001",
"01010001",
"00000110",
"00000000",
"01110001",
"10101001",
"00111010",
"01111110",
"10000101",
"11010100",
"01101100",
"10111010",
"00100010",
"11100010",
"11100111",
"11101100",
"00110100",
"10110111",
"10011001",
"10100000",
"10001111",
"00101000",
"00011100",
"00010101"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;