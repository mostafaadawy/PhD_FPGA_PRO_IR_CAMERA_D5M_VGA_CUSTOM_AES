LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom415 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom415 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom415 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"10001110",
"00101010",
"11110111",
"00011000",
"11000111",
"11001000",
"00101001",
"10111001",
"10111100",
"10110111",
"01010011",
"01111101",
"10110110",
"01001010",
"01000110",
"00111000",
"01101100",
"00010101",
"10001100",
"10000000",
"00001001",
"10010110",
"00011001",
"01101011",
"00001110",
"01101001",
"10001001",
"11010000",
"10010101",
"01110010",
"11110001",
"10010011",
"11001110",
"01010010",
"10000110",
"11111001",
"01011000",
"10110001",
"11110110",
"01001111",
"10010010",
"00100111",
"00110100",
"10011010",
"11111011",
"00111001",
"00111100",
"00001000",
"01100111",
"11101001",
"11010101",
"11110010",
"01100110",
"10101011",
"00010110",
"11001111",
"10111010",
"10100011",
"01111010",
"11100010",
"11101011",
"01111110",
"01001000",
"10010111",
"00011011",
"00101011",
"11010111",
"00100001",
"10011001",
"11100011",
"11110011",
"10001011",
"01001100",
"11111000",
"10011100",
"11011100",
"01101000",
"10100010",
"10101001",
"11000110",
"01110101",
"00000110",
"10011011",
"10100110",
"00100011",
"01101110",
"10101010",
"10011000",
"10011111",
"11101110",
"01001101",
"10111110",
"01001110",
"10101111",
"10101110",
"11000010",
"10110100",
"00110011",
"00000011",
"00110000",
"01000100",
"00001011",
"01011010",
"00101101",
"11001001",
"11000000",
"10000011",
"00111111",
"01100101",
"11101010",
"11011001",
"01010101",
"01010111",
"10111011",
"11101101",
"00001101",
"01100001",
"11001011",
"11101111",
"10110000",
"11000001",
"11000100",
"01000101",
"10100000",
"10001111",
"00100010",
"10010100",
"01011100",
"01111011",
"00010000",
"00111101",
"00001100",
"01000111",
"11011101",
"01011011",
"00011010",
"01000010",
"10010001",
"00011110",
"10111101",
"01000001",
"00011101",
"01001001",
"01011110",
"00010111",
"01110001",
"11110100",
"11010100",
"11001100",
"00101110",
"11111110",
"10111000",
"11011110",
"01101111",
"11100110",
"11111100",
"11100001",
"11111010",
"01100100",
"11001101",
"11010011",
"01000000",
"00001010",
"10101100",
"11010001",
"10100001",
"00011111",
"00000111",
"10000001",
"11011111",
"01000011",
"11101100",
"10000111",
"10101101",
"11100101",
"10100111",
"10011110",
"11010110",
"01111111",
"11011010",
"10100101",
"10101000",
"01110100",
"01101010",
"10001101",
"01011001",
"11110101",
"11111101",
"00000101",
"00010100",
"10000101",
"00000100",
"10110011",
"01110011",
"10001000",
"10100100",
"01001011",
"00010001",
"00110001",
"01011111",
"11001010",
"00010010",
"11110000",
"01010001",
"00110101",
"01011101",
"10011101",
"01100000",
"00100110",
"00111010",
"00110110",
"10000100",
"10110010",
"10110101",
"00010011",
"10010000",
"00101111",
"00111011",
"00000010",
"01010110",
"11000101",
"10000010",
"00111110",
"11011000",
"01111000",
"01010000",
"01111001",
"00101100",
"01101101",
"00101000",
"00100100",
"00011100",
"01010100",
"01110110",
"01100010",
"11100111",
"00110111",
"10001010",
"00100101",
"11100100",
"11101000",
"00000000",
"00110010",
"10111111",
"11010010",
"00001111",
"01110000",
"11011011",
"11100000",
"11111111",
"01110111",
"00000001",
"11000011",
"00100000"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;