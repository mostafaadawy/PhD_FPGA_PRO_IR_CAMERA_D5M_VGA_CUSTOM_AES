LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom319 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom319 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom319 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"10111000",
"00001110",
"11011010",
"11011111",
"11010101",
"11001100",
"10111111",
"11111001",
"01101001",
"00101110",
"01101100",
"10100100",
"11100000",
"10010000",
"00001101",
"00110010",
"01111010",
"10110001",
"01100110",
"01100010",
"10010001",
"10111001",
"10110000",
"11010111",
"10000000",
"11101010",
"11110110",
"01011000",
"10011010",
"11011000",
"01010100",
"11110101",
"11001011",
"11100100",
"11101111",
"01000110",
"01011110",
"11101101",
"10110101",
"10101000",
"11100011",
"11110000",
"00011010",
"10000011",
"01011010",
"01011100",
"11011110",
"01011111",
"01101101",
"00110100",
"10010010",
"00101101",
"11110011",
"11100101",
"10101001",
"01001101",
"10101010",
"01100111",
"10011111",
"01001011",
"10111110",
"11111011",
"11111000",
"01110011",
"00101000",
"11000111",
"00110111",
"10000101",
"10100000",
"10000100",
"00100101",
"01000101",
"11110001",
"01111001",
"11111101",
"00000111",
"00100100",
"00101111",
"00001000",
"11100001",
"11010010",
"10001000",
"01110111",
"11001001",
"11111110",
"01010101",
"10001011",
"10000110",
"00010011",
"01100100",
"10101011",
"10100011",
"11111100",
"01011001",
"11101001",
"00001001",
"01111101",
"11101110",
"00110000",
"00011110",
"10011100",
"00000100",
"10011011",
"11100110",
"00010000",
"10011101",
"01111111",
"10010101",
"00100000",
"00011000",
"01010010",
"10001001",
"01110100",
"11001101",
"11010011",
"00100001",
"00110101",
"01011011",
"01001001",
"11011011",
"00100011",
"10111101",
"10001101",
"00010010",
"01111011",
"10010011",
"11111010",
"00110011",
"01101011",
"10010111",
"11000110",
"11111111",
"01100101",
"10110011",
"00011101",
"00001010",
"01000100",
"11110100",
"11010110",
"00101001",
"11000100",
"01001110",
"00010100",
"00010101",
"01110000",
"10100010",
"01111110",
"01100001",
"01101110",
"11000001",
"00101100",
"11101100",
"01010001",
"01010110",
"10010100",
"10110010",
"00010001",
"01011101",
"10000010",
"10000001",
"01110110",
"10111010",
"10111011",
"11100111",
"10010110",
"10110110",
"00111101",
"00100110",
"00110110",
"01101000",
"10101101",
"10011001",
"01111000",
"10110111",
"00010111",
"01001010",
"11000101",
"00000000",
"00001111",
"10011110",
"10110100",
"11001110",
"01010011",
"00000011",
"01010111",
"10000111",
"10101100",
"10101110",
"00101010",
"11101011",
"01110010",
"01010000",
"00000010",
"00001011",
"00111000",
"10011000",
"10100101",
"00110001",
"11001010",
"00111110",
"11011101",
"01000001",
"11001000",
"01101010",
"11010000",
"10100110",
"00011111",
"11000000",
"10100001",
"11010100",
"10001110",
"11001111",
"01001000",
"00100111",
"00111001",
"11110111",
"01001100",
"00011001",
"11000010",
"11110010",
"10001010",
"11000011",
"10101111",
"01110101",
"00010110",
"01000111",
"10111100",
"11010001",
"01100000",
"11011100",
"00111011",
"00000001",
"01000010",
"10100111",
"00011100",
"00000110",
"00101011",
"01001111",
"00100010",
"11101000",
"00111111",
"11100010",
"01000011",
"00111010",
"00001100",
"10001100",
"01000000",
"01110001",
"10001111",
"11011001",
"01101111",
"00111100",
"00011011",
"00000101"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
