LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom301 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom301 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom301 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type :=(
"01100011",
"01111100",
"01011111",
"10110100",
"01111101",
"11010001",
"10001000",
"01001000",
"11011111",
"10000101",
"00111010",
"10100010",
"10010110",
"11110101",
"01000101",
"00001101",
"10001110",
"01100100",
"10100011",
"01001111",
"11001111",
"00101111",
"00110000",
"11101110",
"00101010",
"11000010",
"00101000",
"00011100",
"01110000",
"11111110",
"01010100",
"00000011",
"00100110",
"01000011",
"01010011",
"10011110",
"10110000",
"00111000",
"01110101",
"00110101",
"10000110",
"10000011",
"11110110",
"11011110",
"11001010",
"10010100",
"10100101",
"10111101",
"11000111",
"11010111",
"10110011",
"10111100",
"11000110",
"01011010",
"11011100",
"00010000",
"11101010",
"11100111",
"10101101",
"10001111",
"11111000",
"10001001",
"11100000",
"01111010",
"01110010",
"01001001",
"11000000",
"10000100",
"11001000",
"01110001",
"00101110",
"00011000",
"00111001",
"10011111",
"11001110",
"00011111",
"11011011",
"11100101",
"11111011",
"11010110",
"00100010",
"11001100",
"00010011",
"11110000",
"10101001",
"00001011",
"00001110",
"00101101",
"10110111",
"10010000",
"00101011",
"00000101",
"00000000",
"01100010",
"00001100",
"01110100",
"10000010",
"11101101",
"10001010",
"01011110",
"10111000",
"00010101",
"10001100",
"00110100",
"00000010",
"01010001",
"01001100",
"10100001",
"00001111",
"00110011",
"01101001",
"01110111",
"00010100",
"00101001",
"00100001",
"01010111",
"00000100",
"10001011",
"10100110",
"11101100",
"00011101",
"10100000",
"00010110",
"11100001",
"00010001",
"00001000",
"11101111",
"01101011",
"11101011",
"10111001",
"11000101",
"01111111",
"10110010",
"10101000",
"00100011",
"10011000",
"10110110",
"00110110",
"01101010",
"11011101",
"01110110",
"11100010",
"01101101",
"10111011",
"01001110",
"10111111",
"10101110",
"10000111",
"00000110",
"01010010",
"01011101",
"10101011",
"00111111",
"11000100",
"00100000",
"11111010",
"10011100",
"01111000",
"00001010",
"00111011",
"11000011",
"00101100",
"00000111",
"11100110",
"11101000",
"10101010",
"00011001",
"01111110",
"10110101",
"01110011",
"11100100",
"00000001",
"11010101",
"00011011",
"11110111",
"01101100",
"00001001",
"01101111",
"10011010",
"10011011",
"01000111",
"11110010",
"01010000",
"10101100",
"01100001",
"01001101",
"11100011",
"10101111",
"11010100",
"11111111",
"01011011",
"01000100",
"10010011",
"00011010",
"00100100",
"10100111",
"10010111",
"00111110",
"11111101",
"01101000",
"00111101",
"01001010",
"01011000",
"10011101",
"00100111",
"11111100",
"01111011",
"10010010",
"01100000",
"11010010",
"11001001",
"00011110",
"11110100",
"11110011",
"10110001",
"00111100",
"01010101",
"11010011",
"01001011",
"00110111",
"01100110",
"10010101",
"11011010",
"11001101",
"11011000",
"01101110",
"01000110",
"11000001",
"01000010",
"01000000",
"01111001",
"01000001",
"11010000",
"11110001",
"00010111",
"00110010",
"10000001",
"10111110",
"10100100",
"01010110",
"01011100",
"10000000",
"00110001",
"11111001",
"11011001",
"00010010",
"10010001",
"10001101",
"11101001",
"01011001",
"01100101",
"11001011",
"00100101",
"10111010",
"01100111",
"10011001"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
