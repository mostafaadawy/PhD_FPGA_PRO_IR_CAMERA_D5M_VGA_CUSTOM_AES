LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom369 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom369 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom369 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"00000110",
"11011010",
"11010001",
"10111000",
"10111111",
"10101110",
"00111010",
"10010100",
"01100100",
"00110101",
"00001101",
"01110001",
"10000101",
"11010101",
"11001111",
"10111101",
"01110010",
"01110100",
"00001010",
"10101111",
"10100010",
"10010010",
"01010100",
"10011101",
"01101010",
"10000010",
"11111010",
"01010001",
"11010010",
"01000011",
"11011111",
"00110000",
"00001100",
"01110111",
"11101011",
"01011110",
"00000010",
"11000001",
"00111101",
"10101010",
"00000101",
"01111010",
"01101001",
"11000011",
"10011011",
"10001011",
"11111000",
"00010010",
"11110110",
"00101001",
"11100111",
"01101110",
"10010011",
"01100001",
"01000101",
"01111111",
"10010000",
"11110010",
"10111011",
"11001000",
"10011001",
"11011000",
"11010111",
"11110101",
"11001010",
"11011001",
"11010100",
"10000110",
"10000011",
"01001001",
"11001101",
"00110111",
"11111101",
"11011011",
"00111001",
"01011111",
"00110010",
"00111000",
"10100110",
"01010111",
"01101101",
"10110011",
"01010000",
"11101001",
"11101111",
"00110100",
"01100110",
"00101110",
"00110011",
"01111110",
"00011111",
"10100111",
"00010111",
"00101011",
"01000100",
"00010001",
"00110001",
"10101101",
"10101001",
"01101111",
"01000110",
"01100101",
"00100001",
"10110001",
"00001111",
"11101000",
"00011011",
"01110110",
"01100010",
"11000100",
"01110000",
"00111011",
"10000111",
"01010011",
"10011010",
"11000110",
"01000001",
"11111100",
"11100101",
"00001001",
"10110110",
"00100100",
"00011110",
"00100111",
"10111110",
"01101000",
"11010011",
"11010110",
"00101000",
"01011100",
"10110111",
"11101101",
"00111110",
"10100000",
"01010010",
"11111110",
"01111011",
"10111010",
"00010011",
"10100001",
"10011100",
"11111001",
"11011110",
"11000010",
"10100011",
"00011000",
"00101100",
"10001100",
"00111111",
"00100110",
"01001110",
"00010110",
"01111101",
"11100010",
"11001011",
"11000111",
"11001110",
"00000000",
"10000001",
"11110111",
"01111001",
"10110010",
"10001110",
"10010101",
"11100001",
"00010100",
"00010000",
"10011110",
"11001100",
"11110011",
"00100101",
"10000100",
"00100010",
"01100111",
"00001011",
"01001101",
"00101111",
"10000000",
"01001011",
"01110101",
"00000111",
"00100011",
"01011101",
"11000101",
"00000001",
"00101101",
"01011001",
"00011010",
"01000111",
"00001110",
"11110000",
"00001000",
"10110000",
"11101110",
"01001010",
"10111001",
"00000100",
"11011100",
"11101100",
"11001001",
"10001111",
"10101000",
"11110001",
"00010101",
"10001010",
"01110011",
"01000010",
"00011001",
"11100000",
"10110100",
"01010101",
"01001000",
"01001100",
"10001000",
"10110101",
"01111000",
"00000011",
"00011100",
"11100011",
"11110100",
"01011010",
"10010110",
"11101010",
"10100100",
"01001111",
"00110110",
"11111011",
"11111111",
"10010001",
"01101100",
"10011111",
"11000000",
"01011011",
"01011000",
"10011000",
"10010111",
"10101100",
"01101011",
"00100000",
"01000000",
"10111100",
"00111100",
"10001001",
"01100000",
"00101010",
"10100101",
"11011101",
"00011101",
"10101011",
"11100100",
"10001101",
"11010000",
"11100110",
"01010110"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
