LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom391 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom391 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom391 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"00001010",
"11010010",
"00110001",
"00001100",
"10111011",
"10010011",
"01001010",
"00110011",
"11010100",
"10001011",
"11101001",
"10111111",
"00011011",
"01000110",
"00010001",
"11000100",
"01001011",
"00010010",
"01011110",
"00101000",
"00010111",
"01101100",
"11000000",
"11001010",
"00001101",
"10101100",
"10111001",
"00111011",
"11110001",
"01000001",
"10111100",
"01111101",
"01010110",
"11100000",
"10010001",
"00101111",
"00111101",
"00010000",
"11111101",
"00000011",
"11000110",
"00000100",
"01011001",
"11011001",
"00000010",
"00100110",
"10110010",
"10000111",
"10110111",
"01000101",
"01010100",
"10110011",
"10000100",
"01010101",
"11101000",
"01100110",
"01001111",
"01011010",
"11001100",
"10101111",
"10010100",
"10100101",
"10001100",
"00100001",
"10001010",
"01100100",
"11111001",
"01011011",
"01000100",
"11011000",
"00011010",
"01101111",
"10100011",
"10011111",
"10101010",
"01110100",
"00111100",
"10011100",
"00101100",
"10011011",
"10110101",
"00111111",
"01010111",
"11000101",
"11010000",
"01110011",
"10011000",
"01110001",
"00111110",
"10100100",
"00110101",
"10000110",
"00100111",
"01101000",
"01101101",
"11110011",
"11110111",
"10010110",
"00001001",
"10100110",
"01110000",
"01011100",
"11111000",
"11110110",
"11101101",
"11111110",
"01110110",
"01100000",
"01111000",
"00011100",
"01000000",
"11100100",
"00000111",
"10010000",
"01110101",
"11011111",
"00011001",
"10110001",
"01010010",
"10110100",
"00000101",
"01000011",
"01111110",
"11111010",
"00000000",
"00101110",
"01110010",
"01011000",
"01000010",
"00010101",
"10010111",
"00011000",
"00000110",
"11101011",
"11001000",
"11000001",
"10011001",
"11010001",
"11110000",
"00111000",
"10111110",
"11111111",
"00111001",
"00111010",
"10000011",
"00011110",
"11100101",
"00110010",
"11111011",
"10110110",
"01100001",
"00101101",
"00001110",
"10001101",
"00101010",
"11001110",
"01111010",
"01001100",
"00100010",
"11011101",
"00011111",
"00010011",
"00001000",
"11001111",
"10101011",
"01001110",
"01111001",
"10001001",
"11010110",
"11001001",
"10111010",
"11001011",
"01101011",
"00100000",
"10011110",
"11110010",
"01101010",
"11010101",
"00101011",
"10100010",
"10000000",
"01100010",
"10101110",
"11110100",
"01110111",
"11101111",
"10100111",
"01010011",
"11100110",
"11000111",
"10000010",
"10111101",
"11001101",
"01011101",
"00101001",
"11011010",
"01111111",
"11000011",
"10110000",
"11110101",
"10000001",
"11100001",
"11101010",
"11010011",
"11111100",
"00110000",
"01001000",
"00110110",
"10101001",
"01011111",
"00100100",
"00010110",
"10101101",
"01101110",
"00001111",
"11000010",
"11100010",
"01100111",
"11101110",
"00110111",
"11011100",
"01101001",
"00010100",
"11011110",
"10100000",
"11100111",
"01010001",
"01001101",
"10011010",
"01111011",
"10001110",
"11100011",
"11011011",
"10010010",
"10111000",
"01100101",
"11101100",
"01000111",
"00011101",
"00100101",
"10001000",
"10001111",
"01010000",
"10101000",
"10010101",
"10000101",
"00001011",
"11010111",
"01001001",
"10100001",
"00110100",
"10011101",
"00100011",
"00000001"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;