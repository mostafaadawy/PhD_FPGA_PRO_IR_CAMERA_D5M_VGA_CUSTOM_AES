LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom333 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom333 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom333 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"01001101",
"01010111",
"01110100",
"10110001",
"01111001",
"11001010",
"01001001",
"00000100",
"10101011",
"11111100",
"01101110",
"11101111",
"10110111",
"00101101",
"11010111",
"01011001",
"11010000",
"00111001",
"10100110",
"01110111",
"10101100",
"00100110",
"01000100",
"01010000",
"00100101",
"01111111",
"00001001",
"00010110",
"11100101",
"01001100",
"10011000",
"10111000",
"11011111",
"11001101",
"10111010",
"10110100",
"01001110",
"10001110",
"10000001",
"10111011",
"11001000",
"10001101",
"10000100",
"01010110",
"01100000",
"01010100",
"11110000",
"11100111",
"01011011",
"01110101",
"11100001",
"01010101",
"11001100",
"00000011",
"11110111",
"01100001",
"11011001",
"00110010",
"00100000",
"01110010",
"11110100",
"01101111",
"10011110",
"01100111",
"00101111",
"01110011",
"10011100",
"10100000",
"10010101",
"10010011",
"00101110",
"10110010",
"10001000",
"10100011",
"11110101",
"01101101",
"00110100",
"11101001",
"00010010",
"11111110",
"10101110",
"00011111",
"10110110",
"10101111",
"10110101",
"10001011",
"00110001",
"01000011",
"11111001",
"10001010",
"11100010",
"11101101",
"11111000",
"01110001",
"00001011",
"00100010",
"00100001",
"11010101",
"11011110",
"00111000",
"11001001",
"00000111",
"10000011",
"11000111",
"01111000",
"10100100",
"00010101",
"01000001",
"11110010",
"11010001",
"00101001",
"10110000",
"01100010",
"10111100",
"00111110",
"01100110",
"11001011",
"01110000",
"11000010",
"10010001",
"11101011",
"11010100",
"10101000",
"11000110",
"11000100",
"11011010",
"00111100",
"00110101",
"11000000",
"10100001",
"11100100",
"10000010",
"01101011",
"00000000",
"00111101",
"01000111",
"00100011",
"11110011",
"10111001",
"11110001",
"00011011",
"10011011",
"01100100",
"00000110",
"00101010",
"11101100",
"10010110",
"11101000",
"10100010",
"00001110",
"00101000",
"01010011",
"11000101",
"00001100",
"01101001",
"01000101",
"10000111",
"10011111",
"01111010",
"11111111",
"10101101",
"01011100",
"10000101",
"00110000",
"01011101",
"01001000",
"10001001",
"01111110",
"00000101",
"00011000",
"00001000",
"10101010",
"00010111",
"10010100",
"01001010",
"00001101",
"11010010",
"10111110",
"10001111",
"11111011",
"10010111",
"01111101",
"00000010",
"01111011",
"00100100",
"11000001",
"00001111",
"11100000",
"01101010",
"01001111",
"11110110",
"00011110",
"11000011",
"01011110",
"01000010",
"01010010",
"10011001",
"01011010",
"00011100",
"00110011",
"11001110",
"11111101",
"00110110",
"10101001",
"01010001",
"11011101",
"00010011",
"11011011",
"10010000",
"10011101",
"11101110",
"01101000",
"10000000",
"10100111",
"01011000",
"00010100",
"11010011",
"00101100",
"00001010",
"11011100",
"00111010",
"01001011",
"01000110",
"10010010",
"00101011",
"00000001",
"11100011",
"10100101",
"10001100",
"11100110",
"01101100",
"10011010",
"01000000",
"10111101",
"00110111",
"11111010",
"11101010",
"00111111",
"10110011",
"11001111",
"00011010",
"11010110",
"10000110",
"01110110",
"00011001",
"00011101",
"00100111",
"00111011",
"00010000",
"01100101",
"00010001",
"01011111",
"10111111",
"11011000"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
