LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY sbox_rom351 IS
   PORT( 
      rom_in  : IN     std_logic_vector (0 TO 7);
      clk     : IN     std_logic;
      rom_out : OUT    std_logic_vector (0 TO 7)
   );

-- Declarations

END sbox_rom351 ;

-- hds interface_end
ARCHITECTURE rtl OF sbox_rom351 IS
Type rom_type is array (0 to 255) of std_logic_vector(0 to 7);
constant rom : rom_type := (
"01100011",
"01111100",
"10101010",
"11101101",
"11000001",
"11100110",
"00100100",
"10001000",
"00110010",
"00111010",
"10100001",
"00111111",
"10000110",
"00110011",
"10010110",
"01100100",
"11001011",
"11100101",
"11001111",
"00010100",
"01000100",
"01000101",
"00001011",
"10101100",
"11010111",
"00111100",
"01001011",
"01010100",
"11011111",
"10101000",
"10100110",
"10000000",
"00110111",
"10111001",
"00100000",
"10100101",
"01110011",
"10111100",
"11011000",
"01011110",
"11110000",
"00011101",
"01110000",
"10101001",
"00010001",
"00001010",
"10000100",
"00101101",
"01111111",
"10100010",
"10001010",
"01100101",
"00110001",
"01001110",
"11111000",
"10011001",
"01111011",
"11011001",
"11000000",
"00001001",
"10000001",
"00101001",
"10010010",
"11111010",
"00001111",
"11101011",
"01001000",
"01101001",
"11000010",
"01000001",
"00000000",
"11011110",
"01101011",
"10111000",
"10001100",
"10001110",
"10111110",
"10111010",
"11111101",
"01001101",
"11101100",
"10111111",
"01011100",
"10100111",
"11101010",
"10011110",
"01000000",
"11001100",
"00011100",
"11001010",
"10010001",
"01100010",
"11010110",
"11000100",
"00000010",
"01111000",
"00101011",
"00110101",
"11000101",
"10101110",
"10010111",
"00100001",
"00100110",
"10000010",
"01001010",
"11110011",
"11110101",
"00110110",
"11101000",
"11111110",
"00011110",
"01010010",
"01101111",
"01011001",
"00111110",
"00111011",
"10110010",
"00000011",
"00010000",
"10111011",
"00010010",
"00101110",
"01000110",
"10110110",
"10011011",
"00100101",
"11101001",
"00100111",
"01010101",
"10100000",
"01100001",
"00110000",
"10110000",
"10011000",
"01100110",
"11011010",
"10110011",
"11010000",
"00110100",
"01011000",
"10010100",
"10101011",
"11111011",
"01110010",
"01100111",
"11101111",
"11001000",
"01110101",
"11010010",
"00101111",
"11010011",
"00010111",
"10001101",
"11010100",
"11001001",
"11001110",
"00101100",
"11100111",
"01110100",
"01000011",
"10100100",
"11110100",
"00001101",
"01010001",
"11111100",
"10100011",
"00000001",
"11100010",
"11100001",
"11000011",
"11011011",
"11010001",
"10110100",
"01101000",
"11110010",
"01011101",
"11011100",
"11110111",
"10110111",
"00010110",
"00011010",
"00111001",
"11100011",
"01101100",
"11111111",
"00111101",
"11110110",
"00010011",
"10010101",
"01010000",
"11101110",
"01011010",
"01000111",
"00101010",
"00001110",
"00011011",
"01110110",
"10011010",
"10000101",
"01010111",
"01011111",
"00001000",
"01000010",
"10110101",
"10000111",
"10010000",
"10010011",
"01111101",
"10110001",
"01111001",
"01101101",
"01010110",
"00101000",
"10011111",
"10001111",
"10101111",
"11100000",
"00011001",
"10101101",
"11010101",
"11011101",
"11000111",
"10111101",
"01110001",
"00100011",
"01101010",
"00111000",
"00001100",
"10001011",
"01110111",
"01001111",
"01111010",
"11001101",
"01111110",
"00010101",
"00000100",
"10011100",
"00011000",
"01001001",
"11100100",
"10011101",
"00000101",
"10000011",
"01010011",
"11110001",
"01011011",
"10001001",
"11000110",
"00011111",
"11111001",
"00000110",
"00100010",
"01100000",
"01101110",
"00000111",
"01001100"
);
BEGIN
process (clk)
variable addr_int: integer range 0 to 255;
begin
  if (rising_edge (clk))then
	addr_int := conv_integer(unsigned(rom_in));
	rom_out <= rom(addr_int);
  end if;
end process;
END rtl;
